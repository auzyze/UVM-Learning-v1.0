/////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////

`ifndef GUARD_CONFIGURATION
`define GUARD_CONFIGURATION

/////////////////////////////////////////////////////////////
// CONFIGURATION FOR SYNC FIFO
/////////////////////////////////////////////////////////////


class my_config extends uvm_object;

`uvm_object_utils(my_config)

bit [3:0]   afull_wtrline;
bit [3:0]   aempt_wtrline;

function new (string name = "");
  super.new(name);
endfunction


endclass :my_config

`endif
