///////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////
///////////  ////////////        //////////////////////////////////
//////////  ///////////////  //////////////////////////////////////
/////////  ///////////////  ///////////////////////////////////////
////////  ///////////////  ////////////////////////////////////////
///////  ///////////////  /////////////////////////////////////////
//////        //////     //////////////////////////////////////////
///////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////


`ifndef GUARD_ENV
`define GUARD_ENV


class environment extends uvm_env;
`uvm_component_utils(environment)

function new(string name, uvm_component parent = null);
  super.new(name, parent);
endfunction


virtual function void build();
  super.build();
  
  uvm_report_info(get_full_name(),"START OF BUILD",UVM_LOW);
  
  uvm_report_info(get_full_name(),"END OF BUILD",UVM_LOW);
    
endfunction


virtual function void connect();
  super.connect();
  
  uvm_report_info(get_full_name(),"START OF CONNECT",UVM_LOW);
  
  uvm_report_info(get_full_name(),"END OF CONNECT",UVM_LOW);
  
endfunction


endclass

`endif

`endif
