//transactions are the basic data objects that are passed between components
