///////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////
///////////  ////////////        //////////////////////////////////
//////////  ///////////////  //////////////////////////////////////
/////////  ///////////////  ///////////////////////////////////////
////////  ///////////////  ////////////////////////////////////////
///////  ///////////////  /////////////////////////////////////////
//////        //////     //////////////////////////////////////////
///////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////

`ifndef GUARD_CONFIGURATION
`define GUARD_CONFIGURATION

/////////////////////////////////////////////////////////////
// CONFIGURATION FOR ASYNC FIFO
/////////////////////////////////////////////////////////////


class my_config extends uvm_object;

`uvm_object_utils(my_config)


/////////////////////////////////////////////////////////////
// virtual interface
//

/////////////////////////////////////////////////////////////
//Using a virtual interface as a reference or handle to the interface instance, 
//the testbench can access the tasks, functions, ports, and internal variables of the
//SystemVerilog interface. ---- from "COOKBOOK" p83


/////////////////////////////////////////////////////////////
//The example of using virtual interface in a Driver. 
//-----see "COOKBOOK" p86


//Declare All the interfaces which are required in this verification environment.

//Used by other verification components like "drive" "moniter" to access physical
//interface in top module using configuration class object ???

virtual fifo_interface.WR wr_intf;
virtual fifo_interface.RD rd_intf;

bit [3:0]   afull_wtrline;
bit [3:0]   aempt_wtrline;


/////////////////////////////////////////////////////////////
//?????????????????????
//what does "this" indicate ??
//why return a "t" ??
//how does the "update" happen ??
//
virtual function uvm_object_create(string name = "");
  my_config t = new();
  
  t.afull_wtrline = this.afull_wtrline;
  t.aempt_wtrline = this.aempt_wtrline;
  t.wr_intf = this.wr_intf;
  t.rd_intf = this.rd_intf;

return t;
endfunction;create

//function new (string name = "");
//  super.new(name);
//endfunction


endclass:my_config

`endif
